netcdf aod_obs_2015081000_m {
dimensions:
	nobs = 1100 ;
	Observation_Class_maxstrlen = 7 ;
	nchans = 11 ;
	nlocs = 100 ;
	nrecs = 100 ;
	nvars = 11 ;
variables:
	int record_number(nlocs) ;
	int chaninfoidx(nchans) ;
	double frequency(nchans) ;
	double polarization(nchans) ;
	double wavenumber(nchans) ;
	double error_variance(nchans) ;
	int use_flag(nchans) ;
	int sensor_chan(nchans) ;
	int satinfo_chan(nchans) ;
	double latitude(nlocs) ;
	double longitude(nlocs) ;
	double time(nlocs) ;
	double Sol_Zenith_Angle(nlocs) ;
	double Sol_Azimuth_Angle(nlocs) ;
	double aerosol_optical_depth_1_(nlocs) ;
	double aerosol_optical_depth_2_(nlocs) ;
	double aerosol_optical_depth_3_(nlocs) ;
	double aerosol_optical_depth_4_(nlocs) ;
	double aerosol_optical_depth_5_(nlocs) ;
	double aerosol_optical_depth_6_(nlocs) ;
	double aerosol_optical_depth_7_(nlocs) ;
	double aerosol_optical_depth_8_(nlocs) ;
	double aerosol_optical_depth_9_(nlocs) ;
	double aerosol_optical_depth_10_(nlocs) ;
	double aerosol_optical_depth_11_(nlocs) ;
	double aerosol_optical_depth_err_1_(nlocs) ;
	double aerosol_optical_depth_err_2_(nlocs) ;
	double aerosol_optical_depth_err_3_(nlocs) ;
	double aerosol_optical_depth_err_4_(nlocs) ;
	double aerosol_optical_depth_err_5_(nlocs) ;
	double aerosol_optical_depth_err_6_(nlocs) ;
	double aerosol_optical_depth_err_7_(nlocs) ;
	double aerosol_optical_depth_err_8_(nlocs) ;
	double aerosol_optical_depth_err_9_(nlocs) ;
	double aerosol_optical_depth_err_10_(nlocs) ;
	double aerosol_optical_depth_err_11_(nlocs) ;
	double aerosol_optical_depth_qc_1_(nlocs) ;
	double aerosol_optical_depth_qc_2_(nlocs) ;
	double aerosol_optical_depth_qc_3_(nlocs) ;
	double aerosol_optical_depth_qc_4_(nlocs) ;
	double aerosol_optical_depth_qc_5_(nlocs) ;
	double aerosol_optical_depth_qc_6_(nlocs) ;
	double aerosol_optical_depth_qc_7_(nlocs) ;
	double aerosol_optical_depth_qc_8_(nlocs) ;
	double aerosol_optical_depth_qc_9_(nlocs) ;
	double aerosol_optical_depth_qc_10_(nlocs) ;
	double aerosol_optical_depth_qc_11_(nlocs) ;
	double obs_minus_forecast_unadjusted_1_(nlocs) ;
	double obs_minus_forecast_unadjusted_2_(nlocs) ;
	double obs_minus_forecast_unadjusted_3_(nlocs) ;
	double obs_minus_forecast_unadjusted_4_(nlocs) ;
	double obs_minus_forecast_unadjusted_5_(nlocs) ;
	double obs_minus_forecast_unadjusted_6_(nlocs) ;
	double obs_minus_forecast_unadjusted_7_(nlocs) ;
	double obs_minus_forecast_unadjusted_8_(nlocs) ;
	double obs_minus_forecast_unadjusted_9_(nlocs) ;
	double obs_minus_forecast_unadjusted_10_(nlocs) ;
	double obs_minus_forecast_unadjusted_11_(nlocs) ;
	double surface_air_pressure_1_(nlocs) ;
	double surface_air_pressure_2_(nlocs) ;
	double surface_air_pressure_3_(nlocs) ;
	double surface_air_pressure_4_(nlocs) ;
	double surface_air_pressure_5_(nlocs) ;
	double surface_air_pressure_6_(nlocs) ;
	double surface_air_pressure_7_(nlocs) ;
	double surface_air_pressure_8_(nlocs) ;
	double surface_air_pressure_9_(nlocs) ;
	double surface_air_pressure_10_(nlocs) ;
	double surface_air_pressure_11_(nlocs) ;

// global attributes:
		:Satellite_Sensor = "v.viirs-m_npp" ;
		:Satellite = "viirs" ;
		:Observation_type = "viirs_aod" ;
		:Outer_Loop_Iteration = 1 ;
		:Number_of_channels = 11 ;
		:date_time = 2018041500 ;
		:ireal_aoddiag = 6 ;
		:ipchan_aoddiag = 4 ;
		:ioff0 = 0 ;
		:history = "Tue Mar 13 13:15:48 2018: ncks -F -d nobs,1,1100 diag_viirs_ges.2015081000_dbl.nc4 diag_viirs_ges.2015081000_dbl_subset.nc4" ;
		:NCO = "4.6.6" ;
data:

 record_number = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100 ;

 chaninfoidx = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11 ;

 frequency = 730328.125, 676117.375, 617006.625, 544471.4375, 446615.28125, 
    402298.40625, 348017.53125, 242116.875, 217983.125, 187270.75, 
    132836.203125 ;

 polarization = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wavenumber = 24361.125, 22552.84765625, 20581.125, 18161.61328125, 
    14897.482421875, 13419.23046875, 11608.615234375, 8076.14990234375, 
    7271.134765625, 6246.6796875, 4430.93896484375 ;

 error_variance = 0.0500000007450581, 0.0500000007450581, 0.0500000007450581, 
    0.0500000007450581, 0.0500000007450581, 0.0500000007450581, 
    0.0500000007450581, 0.0500000007450581, 0.0500000007450581, 
    0.0500000007450581, 0.0500000007450581 ;

 use_flag = -1, -1, -1, 1, -1, -1, -1, -1, -1, -1, -1 ;

 sensor_chan = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11 ;

 satinfo_chan = 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51 ;

 latitude = 64.5886535644531, 64.6759872436523, 65.1799163818359, 
    65.1146926879883, 65.3409805297852, 65.2393264770508, 65.8974380493164, 
    65.8558120727539, 66.0940628051758, 66.1785583496094, 66.144401550293, 
    66.9555969238281, 67.1115036010742, 66.9841384887695, 68.0091323852539, 
    67.9401168823242, 67.8942413330078, 68.6528091430664, 68.9857788085938, 
    70.036979675293, 69.9070205688477, 70.3742828369141, 70.5062637329102, 
    76.4745101928711, 76.2386703491211, 75.806022644043, 77.2142562866211, 
    76.8106994628906, 78.2385101318359, 79.0149917602539, 78.8103485107422, 
    79.5588607788086, 79.7070083618164, 65.5009384155273, 65.0460433959961, 
    66.362663269043, 66.35009765625, 67.1916732788086, 67.0661697387695, 
    67.0972900390625, 67.1482086181641, 66.9544830322266, 67.3707733154297, 
    67.0068588256836, 67.0188217163086, 67.8101272583008, 67.8502426147461, 
    68.0246963500977, 67.5010070800781, 67.7971572875977, 67.6376113891602, 
    68.7847213745117, 68.8718338012695, 68.4190902709961, 69.0947799682617, 
    69.6169662475586, 69.662971496582, 69.6843872070312, 70.6279830932617, 
    70.5858993530273, 70.4176177978516, 70.7197418212891, 71.0281982421875, 
    71.6572036743164, 71.5176391601562, 71.7996063232422, 71.8094863891602, 
    71.7812271118164, 71.7633972167969, 72.3242416381836, 72.3352966308594, 
    72.4318084716797, 72.4687118530273, 72.2579879760742, 73.6514663696289, 
    73.9417037963867, 74.3609619140625, 76.4003067016602, 76.9257278442383, 
    79.9178466796875, 79.6632919311523, 80.557991027832, 80.4627380371094, 
    64.4303894042969, 66.1602935791016, 67.3615112304688, 67.3844985961914, 
    66.8545913696289, 67.9791030883789, 67.7731704711914, 67.6170501708984, 
    67.8195266723633, 71.8471298217773, 71.9156188964844, 72.8270797729492, 
    72.463623046875, 72.8214874267578, 73.0835723876953, 73.2235336303711, 
    73.4597930908203 ;

 longitude = 51.4124717712402, 51.9743499755859, 48.9114112854004, 
    49.963508605957, 52.3498001098633, 54.6642189025879, 47.6314010620117, 
    49.2311897277832, 52.2236404418945, 54.5701217651367, 55.6933708190918, 
    49.1902885437012, 51.5516014099121, 54.1682510375977, 49.1846084594727, 
    51.1826210021973, 54.1439208984375, 51.4869613647461, 52.9109001159668, 
    50.4959182739258, 52.1353912353516, 51.0901298522949, 52.5974388122559, 
    40.7710494995117, 41.613899230957, 53.5627784729004, 39.5261306762695, 
    41.1086807250977, 48.7806701660156, 44.7753295898438, 48.2780609130859, 
    48.653980255127, 50.4320297241211, 56.1118011474609, 78.150390625, 
    72.9782867431641, 74.2277221679688, 56.3336601257324, 58.2549705505371, 
    60.1977005004883, 70.3084564208984, 72.5562210083008, 73.8848724365234, 
    77.4877395629883, 79.7254486083984, 55.9332809448242, 68.5817337036133, 
    71.0502090454102, 72.8478469848633, 74.5447692871094, 77.0992202758789, 
    67.9930419921875, 70.6088562011719, 74.2179565429688, 75.4262084960938, 
    71.2907867431641, 73.1902084350586, 76.0687637329102, 72.9528427124023, 
    74.0945587158203, 77.0968322753906, 79.8847732543945, 81.2661972045898, 
    70.1412582397461, 72.2285766601562, 75.7224197387695, 78.1791534423828, 
    81.4773788452148, 83.1796264648438, 70.3921737670898, 73.5185928344727, 
    75.8486175537109, 79.2280426025391, 81.6354064941406, 74.2146987915039, 
    74.3828506469727, 76.6857223510742, 71.4002532958984, 72.0137634277344, 
    56.4575996398926, 60.2137298583984, 63.2261581420898, 76.9067230224609, 
    99.7358703613281, 110.63215637207, 95.8495101928711, 97.1000518798828, 
    110.432441711426, 94.92578125, 96.7880172729492, 108.584136962891, 
    110.250129699707, 85.9896392822266, 88.1573028564453, 84.202507019043, 
    87.5781021118164, 89.6472396850586, 83.9737167358398, 85.8865966796875, 
    89.5709991455078 ;

 time = -0.816666662693024, -0.816666662693024, -0.816666662693024, 
    -0.816666662693024, -0.833333313465118, -0.833333313465118, 
    -0.816666662693024, -0.816666662693024, -0.833333313465118, 
    -0.833333313465118, -0.833333313465118, -0.816666662693024, 
    -0.833333313465118, -0.833333313465118, -0.833333313465118, 
    -0.833333313465118, -0.833333313465118, -0.833333313465118, 
    -0.833333313465118, -0.833333313465118, -0.833333313465118, 
    -0.833333313465118, -0.833333313465118, -0.833333313465118, 
    -0.833333313465118, -0.850000023841858, -0.833333313465118, 
    -0.833333313465118, -0.850000023841858, -0.850000023841858, 
    -0.850000023841858, -0.850000023841858, -0.850000023841858, 
    -0.833333313465118, -2.51666665077209, -2.51666665077209, 
    -2.51666665077209, -0.833333313465118, -0.833333313465118, 
    -0.833333313465118, -0.850000023841858, -2.51666665077209, 
    -2.51666665077209, -2.51666665077209, -2.51666665077209, 
    -0.833333313465118, -0.850000023841858, -0.850000023841858, 
    -2.51666665077209, -2.51666665077209, -2.51666665077209, 
    -0.850000023841858, -2.51666665077209, -2.51666665077209, 
    -2.51666665077209, -2.51666665077209, -2.51666665077209, 
    -2.51666665077209, -2.51666665077209, -2.51666665077209, 
    -0.883333325386047, -2.53333330154419, -2.53333330154419, 
    -0.850000023841858, -2.51666665077209, -2.51666665077209, 
    -0.883333325386047, -2.53333330154419, -2.53333330154419, 
    -2.51666665077209, -2.51666665077209, -2.51666665077209, 
    -2.53333330154419, -2.53333330154419, -2.51666665077209, 
    -2.53333330154419, -0.883333325386047, -0.850000023841858, 
    -2.53333330154419, -2.53333330154419, -2.53333330154419, 
    -2.53333330154419, -2.53333330154419, -4.19999980926514, 
    -4.21666669845581, -2.53333330154419, -2.53333330154419, 
    -4.21666669845581, -0.899999976158142, -2.53333330154419, 
    -4.21666669845581, -2.56666660308838, -0.883333325386047, 
    -2.53333330154419, -0.883333325386047, -2.53333330154419, 
    -0.883333325386047, -2.53333330154419, -0.883333325386047, 
    -2.53333330154419 ;

 Sol_Zenith_Angle = 76.9599990844727, 77.4599990844727, 74.9000015258789, 
    75.8000030517578, 77.9000015258789, 79.8899993896484, 73.8899993896484, 
    75.2799987792969, 77.9300003051758, 79.9899978637695, 80.9700012207031, 
    75.4100036621094, 77.5100021362305, 79.7900009155273, 75.5699996948242, 
    77.3300018310547, 79.9499969482422, 77.7300033569336, 79.0599975585938, 
    77.0800018310547, 78.5400009155273, 77.6800003051758, 79.0800018310547, 
    69.0999984741211, 69.8600006103516, 81.0500030517578, 68.0299987792969, 
    69.4700012207031, 77.0100021362305, 73.3199996948242, 76.6399993896484, 
    77.1500015258789, 78.8899993896484, 81.2099990844727, 78.2099990844727, 
    73.9199981689453, 75.0100021362305, 81.75, 83.4300003051758, 
    85.1600036621094, 94.2399978637695, 73.629997253418, 74.8600006103516, 
    77.9800033569336, 79.9499969482422, 81.5299987792969, 92.9000015258789, 
    95.1999969482422, 73.9599990844727, 75.5100021362305, 77.75, 
    92.6500015258789, 72.1600036621094, 75.3199996948242, 76.5100021362305, 
    72.879997253418, 74.5999984741211, 77.1900024414062, 74.5299987792969, 
    75.5599975585938, 101.669998168945, 80.8499984741211, 82.1800003051758, 
    95.5400009155273, 74.0100021362305, 77.25, 103.209999084473, 
    82.5299987792969, 84.0999984741211, 72.4499969482422, 75.3300018310547, 
    77.4800033569336, 80.6100006103516, 82.7900009155273, 76.1999969482422, 
    76.4100036621094, 102.690002441406, 98.25, 74.7200012207031, 
    60.3199996948242, 63.8899993896484, 66.9199981689453, 80.120002746582, 
    74.8399963378906, 84.629997253418, 94.4499969482422, 95.5999984741211, 
    84.620002746582, 117.839996337891, 95.4499969482422, 83.1600036621094, 
    108, 110.769996643066, 88.75, 109.410003662109, 88.3499984741211, 
    114.76000213623, 85.1500015258789, 111.209999084473, 90.5 ;

 Sol_Azimuth_Angle = 3, 1, 3, 1, 1, 3, 1, 1, 3, 1, 1, 1, 3, 3, 0, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 
    1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 0, 0, 1, 0, 1, 0, 0, 1, 1, 1, 1, 0, 0, 3, 
    0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 3, 3, 2, 2, 2, 3, 
    2, 1, 3, 0, 1, 1, 2, 2, 1 ;

 aerosol_optical_depth_1_ = 0.0710000023245811, 0.0489999987185001, 
    0.112000003457069, 0.0750000029802322, 0.0450000017881393, 
    0.0540000014007092, 0.0509999990463257, 0.0529999993741512, 
    0.158999994397163, 0.0549999997019768, 0.028999999165535, 
    0.0850000008940697, 0.108000002801418, 0.158000007271767, 
    0.061999998986721, 0.122000001370907, 0.0520000010728836, 
    0.0869999974966049, 0.0850000008940697, 0.0549999997019768, 
    0.034000001847744, 0.146999999880791, 0.123000003397465, 
    0.0540000014007092, 0.0740000009536743, 0.0309999994933605, 
    0.0370000004768372, 0.0309999994933605, 0.0520000010728836, 
    0.0230000000447035, 0.0390000008046627, 0.0430000014603138, 
    0.0320000015199184, 0.0410000011324883, 0.0769999995827675, 
    0.0379999987781048, 0.0399999991059303, 0.129999995231628, 
    0.0270000007003546, 0.0399999991059303, 0.0399999991059303, 
    0.0729999989271164, 0.0450000017881393, 0.0189999993890524, 
    0.0790000036358833, 0.0689999982714653, 0.063000001013279, 
    0.105999998748302, 0.0670000016689301, 0.0520000010728836, 
    0.00800000037997961, 0.0549999997019768, 0.0149999996647239, 
    0.0329999998211861, 0.0430000014603138, 0.0350000001490116, 
    0.0750000029802322, 0.0219999998807907, 0.0810000002384186, 
    0.0710000023245811, 0.025000000372529, 0.0890000015497208, 
    0.0359999984502792, 0.00400000018998981, 0.0689999982714653, 
    0.115000002086163, 0.00100000004749745, 0.0790000036358833, 
    0.0390000008046627, 0.0209999997168779, 0.0750000029802322, 
    0.0890000015497208, 0.0719999969005585, 0.0450000017881393, 
    0.0379999987781048, 0.034000001847744, 0.0540000014007092, 
    0.0790000036358833, 0.0160000007599592, 0.119999997317791, 
    0.293000012636185, 0.0790000036358833, 0.225999996066093, 
    0.119999997317791, 0.120999999344349, 0.226999998092651, 
    0.26800000667572, 0.0989999994635582, 0.310999989509583, 
    0.221000000834465, 0.138999998569489, 0.20100000500679, 
    0.122000001370907, 0.465999990701675, 0.101999998092651, 
    0.0489999987185001, 0.0570000000298023, 0.028999999165535, 
    0.00899999961256981, 0.0130000002682209 ;

 aerosol_optical_depth_2_ = 0.063000001013279, 0.0469999983906746, 
    0.100000001490116, 0.0719999969005585, 0.0439999997615814, 
    0.0480000004172325, 0.0489999987185001, 0.0509999990463257, 
    0.14300000667572, 0.0529999993741512, 0.0280000008642673, 
    0.0810000002384186, 0.0970000028610229, 0.141000002622604, 
    0.0570000000298023, 0.116999998688698, 0.0500000007450581, 
    0.0799999982118607, 0.0790000036358833, 0.0469999983906746, 
    0.0309999994933605, 0.13400000333786, 0.115000002086163, 
    0.046000000089407, 0.0659999996423721, 0.0280000008642673, 
    0.034000001847744, 0.0270000007003546, 0.0439999997615814, 
    0.0199999995529652, 0.0329999998211861, 0.0370000004768372, 
    0.0280000008642673, 0.0399999991059303, 0.0740000009536743, 
    0.0370000004768372, 0.0379999987781048, 0.123999997973442, 
    0.0260000005364418, 0.0379999987781048, 0.0390000008046627, 
    0.063000001013279, 0.0410000011324883, 0.0179999992251396, 
    0.0759999975562096, 0.0659999996423721, 0.0599999986588955, 
    0.0949999988079071, 0.0570000000298023, 0.0469999983906746, 
    0.00700000021606684, 0.0520000010728836, 0.0140000004321337, 
    0.0299999993294477, 0.0390000008046627, 0.034000001847744, 
    0.0640000030398369, 0.0209999997168779, 0.0689999982714653, 
    0.061999998986721, 0.0240000002086163, 0.0850000008940697, 
    0.034000001847744, 0.00400000018998981, 0.0599999986588955, 
    0.101000003516674, 0.00100000004749745, 0.0689999982714653, 
    0.0379999987781048, 0.0179999992251396, 0.0640000030398369, 
    0.0759999975562096, 0.0649999976158142, 0.0419999994337559, 
    0.0359999984502792, 0.0320000015199184, 0.0489999987185001, 
    0.0769999995827675, 0.0149999996647239, 0.103000000119209, 
    0.261000007390976, 0.068000003695488, 0.195999994874001, 
    0.115000002086163, 0.108000002801418, 0.202999994158745, 
    0.24099999666214, 0.0879999995231628, 0.27700001001358, 
    0.195999994874001, 0.123999997973442, 0.179000005125999, 
    0.116999998688698, 0.419999986886978, 0.0970000028610229, 
    0.0469999983906746, 0.0549999997019768, 0.0260000005364418, 
    0.00800000037997961, 0.0130000002682209 ;

 aerosol_optical_depth_3_ = 0.0549999997019768, 0.0439999997615814, 
    0.0860000029206276, 0.0670000016689301, 0.0410000011324883, 
    0.0410000011324883, 0.046000000089407, 0.0480000004172325, 
    0.123000003397465, 0.0489999987185001, 0.0260000005364418, 
    0.0759999975562096, 0.0829999968409538, 0.122000001370907, 
    0.0500000007450581, 0.108999997377396, 0.046000000089407, 
    0.0710000023245811, 0.0719999969005585, 0.0379999987781048, 
    0.0270000007003546, 0.119999997317791, 0.104000002145767, 
    0.0370000004768372, 0.0570000000298023, 0.0230000000447035, 
    0.0299999993294477, 0.0219999998807907, 0.0359999984502792, 
    0.0160000007599592, 0.0270000007003546, 0.0299999993294477, 
    0.0240000002086163, 0.0370000004768372, 0.0689999982714653, 
    0.034000001847744, 0.0359999984502792, 0.11599999666214, 
    0.0240000002086163, 0.0359999984502792, 0.0359999984502792, 
    0.0520000010728836, 0.0370000004768372, 0.017000000923872, 
    0.0710000023245811, 0.0610000006854534, 0.0560000017285347, 
    0.0820000022649765, 0.046000000089407, 0.0419999994337559, 
    0.00700000021606684, 0.0480000004172325, 0.0130000002682209, 
    0.0270000007003546, 0.0350000001490116, 0.0309999994933605, 
    0.0529999993741512, 0.0199999995529652, 0.0570000000298023, 
    0.0509999990463257, 0.0219999998807907, 0.0790000036358833, 
    0.0320000015199184, 0.00400000018998981, 0.0500000007450581, 
    0.0860000029206276, 0, 0.0579999983310699, 0.0359999984502792, 
    0.0160000007599592, 0.0520000010728836, 0.063000001013279, 
    0.0560000017285347, 0.0379999987781048, 0.034000001847744, 
    0.028999999165535, 0.0439999997615814, 0.0740000009536743, 
    0.0149999996647239, 0.0850000008940697, 0.225999996066093, 
    0.0560000017285347, 0.163000002503395, 0.10700000077486, 
    0.0930000022053719, 0.174999997019768, 0.208000004291534, 
    0.0750000029802322, 0.238000005483627, 0.167999997735023, 
    0.10700000077486, 0.152999997138977, 0.108999997377396, 
    0.365000009536743, 0.0900000035762787, 0.0439999997615814, 
    0.0509999990463257, 0.0219999998807907, 0.00700000021606684, 
    0.0120000001043081 ;

 aerosol_optical_depth_4_ = 0.0209999997168779, 0.017000000923872, 
    0.0784000009298325, 0.0670399963855743, 0.0140000004321337, 
    0.0109999999403954, 0.0189999993890524, 0.0209999997168779, 
    0.119580000638962, 0.0219999998807907, 0.00100000004749745, 
    0.0784000009298325, 0.0741399973630905, 0.118160001933575, 
    0.0199999995529652, 0.122419998049736, 0.0199999995529652, 
    0.0379999987781048, 0.0399999991059303, 0.00700000021606684, 
    0.00100000004749745, 0.0829999968409538, 0.068000003695488, 
    0.00600000005215406, 0.025000000372529, 0, 0.00400000018998981, 0, 
    0.00499999988824129, 0, 0, 0, 0, 0.0109999999403954, 0.0684600025415421, 
    0.00800000037997961, 0.00999999977648258, 0.13094000518322, 0, 
    0.00999999977648258, 0.00999999977648258, 0.017000000923872, 
    0.00899999961256981, 0, 0.0712999999523163, 0.0585200004279613, 
    0.0528399981558323, 0.0469999983906746, 0.0120000001043081, 
    0.0130000002682209, 0, 0.0209999997168779, 0, 0.00100000004749745, 
    0.00700000021606684, 0.00600000005215406, 0.0179999992251396, 0, 
    0.0209999997168779, 0.017000000923872, 0, 0.0826599970459938, 
    0.00600000005215406, 0, 0.0160000007599592, 0.0469999983906746, 0, 
    0.0240000002086163, 0.0109999999403954, 0, 0.017000000923872, 
    0.025000000372529, 0.025000000372529, 0.00999999977648258, 
    0.00899999961256981, 0.00400000018998981, 0.0149999996647239, 
    0.0480000004172325, 0, 0.0439999997615814, 0.165999993681908, 
    0.0209999997168779, 0.104999996721745, 0.119580000638962, 
    0.0840800032019615, 0.180639997124672, 0.187000006437302, 
    0.0656199976801872, 0.210999995470047, 0.170699998736382, 
    0.102540001273155, 0.153659999370575, 0.120999999344349, 
    0.316000014543533, 0.0579999983310699, 0.017000000923872, 
    0.0240000002086163, 0, 0, 0 ;

 aerosol_optical_depth_5_ = 0.0309999994933605, 0.0350000001490116, 
    0.0480000004172325, 0.0540000014007092, 0.0329999998211861, 
    0.0230000000447035, 0.0370000004768372, 0.0379999987781048, 
    0.0689999982714653, 0.0390000008046627, 0.0209999997168779, 
    0.0610000006854534, 0.0469999983906746, 0.068000003695488, 
    0.0299999993294477, 0.0890000015497208, 0.0370000004768372, 
    0.0439999997615814, 0.0469999983906746, 0.0179999992251396, 
    0.0179999992251396, 0.0869999974966049, 0.0689999982714653, 
    0.0160000007599592, 0.0350000001490116, 0.0140000004321337, 
    0.0189999993890524, 0.0109999999403954, 0.0160000007599592, 
    0.00700000021606684, 0.0120000001043081, 0.0130000002682209, 
    0.0140000004321337, 0.0299999993294477, 0.0549999997019768, 
    0.0270000007003546, 0.028999999165535, 0.0939999967813492, 
    0.0189999993890524, 0.0280000008642673, 0.028999999165535, 
    0.025000000372529, 0.0230000000447035, 0.0140000004321337, 
    0.0570000000298023, 0.0489999987185001, 0.0450000017881393, 
    0.0529999993741512, 0.0199999995529652, 0.025000000372529, 
    0.00499999988824129, 0.0359999984502792, 0.00999999977648258, 
    0.0179999992251396, 0.0209999997168779, 0.025000000372529, 
    0.0260000005364418, 0.0160000007599592, 0.0270000007003546, 
    0.0260000005364418, 0.0179999992251396, 0.0640000030398369, 
    0.025000000372529, 0.00300000002607703, 0.025000000372529, 
    0.0500000007450581, 0, 0.0329999998211861, 0.028999999165535, 
    0.00899999961256981, 0.0240000002086163, 0.028999999165535, 
    0.0359999984502792, 0.025000000372529, 0.0260000005364418, 
    0.0209999997168779, 0.0270000007003546, 0.0649999976158142, 
    0.0140000004321337, 0.0430000014603138, 0.143999993801117, 
    0.0270000007003546, 0.0850000008940697, 0.0869999974966049, 
    0.0520000010728836, 0.0979999974370003, 0.116999998688698, 
    0.0419999994337559, 0.13400000333786, 0.0939999967813492, 
    0.0599999986588955, 0.0860000029206276, 0.0890000015497208, 
    0.208000004291534, 0.063000001013279, 0.0350000001490116, 
    0.0410000011324883, 0.0130000002682209, 0.00400000018998981, 
    0.00999999977648258 ;

 aerosol_optical_depth_6_ = 0.025000000372529, 0.0329999998211861, 
    0.0390000008046627, 0.0509999990463257, 0.0309999994933605, 
    0.0189999993890524, 0.034000001847744, 0.0359999984502792, 
    0.0560000017285347, 0.0370000004768372, 0.0189999993890524, 
    0.0579999983310699, 0.0379999987781048, 0.0549999997019768, 
    0.025000000372529, 0.0839999988675117, 0.0350000001490116, 
    0.0370000004768372, 0.0399999991059303, 0.0140000004321337, 
    0.0160000007599592, 0.0799999982118607, 0.0590000003576279, 
    0.0120000001043081, 0.0309999994933605, 0.0120000001043081, 
    0.0160000007599592, 0.00899999961256981, 0.0120000001043081, 
    0.00499999988824129, 0.00899999961256981, 0.00999999977648258, 
    0.0120000001043081, 0.0280000008642673, 0.0520000010728836, 
    0.0260000005364418, 0.0270000007003546, 0.0900000035762787, 
    0.0179999992251396, 0.0270000007003546, 0.0270000007003546, 
    0.0189999993890524, 0.0189999993890524, 0.0130000002682209, 
    0.0540000014007092, 0.0469999983906746, 0.0430000014603138, 
    0.046000000089407, 0.0149999996647239, 0.0199999995529652, 
    0.00499999988824129, 0.0329999998211861, 0.00999999977648258, 
    0.0149999996647239, 0.0179999992251396, 0.0230000000447035, 
    0.0199999995529652, 0.0149999996647239, 0.0209999997168779, 
    0.0209999997168779, 0.0160000007599592, 0.0610000006854534, 
    0.0240000002086163, 0.00300000002607703, 0.0209999997168779, 
    0.0430000014603138, 0, 0.0280000008642673, 0.0270000007003546, 
    0.00700000021606684, 0.0189999993890524, 0.0230000000447035, 
    0.0320000015199184, 0.0219999998807907, 0.0230000000447035, 
    0.0189999993890524, 0.0219999998807907, 0.061999998986721, 
    0.0140000004321337, 0.034000001847744, 0.128000006079674, 
    0.0209999997168779, 0.0689999982714653, 0.0829999968409538, 
    0.0430000014603138, 0.0799999982118607, 0.0949999988079071, 
    0.0350000001490116, 0.109999999403954, 0.0780000016093254, 
    0.0489999987185001, 0.0710000023245811, 0.0839999988675117, 
    0.168999999761581, 0.0549999997019768, 0.0329999998211861, 
    0.0390000008046627, 0.00999999977648258, 0.00300000002607703, 
    0.00899999961256981 ;

 aerosol_optical_depth_7_ = 0.0189999993890524, 0.0299999993294477, 
    0.0299999993294477, 0.0480000004172325, 0.0280000008642673, 
    0.0149999996647239, 0.0320000015199184, 0.0329999998211861, 
    0.0419999994337559, 0.0350000001490116, 0.0179999992251396, 
    0.0540000014007092, 0.028999999165535, 0.0419999994337559, 
    0.0189999993890524, 0.0790000036358833, 0.0320000015199184, 
    0.028999999165535, 0.0320000015199184, 0.00899999961256981, 
    0.0149999996647239, 0.0719999969005585, 0.0469999983906746, 
    0.00800000037997961, 0.0270000007003546, 0.00999999977648258, 
    0.0120000001043081, 0.00700000021606684, 0.00800000037997961, 
    0.00300000002607703, 0.00600000005215406, 0.00600000005215406, 
    0.00999999977648258, 0.0260000005364418, 0.0489999987185001, 
    0.0240000002086163, 0.025000000372529, 0.0839999988675117, 
    0.0160000007599592, 0.025000000372529, 0.025000000372529, 
    0.0140000004321337, 0.0149999996647239, 0.0120000001043081, 
    0.0500000007450581, 0.0430000014603138, 0.0399999991059303, 
    0.0399999991059303, 0.00999999977648258, 0.0149999996647239, 
    0.00499999988824129, 0.0299999993294477, 0.00899999961256981, 
    0.0120000001043081, 0.0140000004321337, 0.0219999998807907, 
    0.0149999996647239, 0.0130000002682209, 0.0149999996647239, 
    0.0149999996647239, 0.0149999996647239, 0.0570000000298023, 
    0.0219999998807907, 0.00300000002607703, 0.0160000007599592, 
    0.0359999984502792, 0, 0.0230000000447035, 0.0240000002086163, 
    0.00600000005215406, 0.0130000002682209, 0.0160000007599592, 
    0.0270000007003546, 0.0179999992251396, 0.0199999995529652, 
    0.017000000923872, 0.017000000923872, 0.0590000003576279, 
    0.0140000004321337, 0.025000000372529, 0.112999998033047, 
    0.0149999996647239, 0.0529999993741512, 0.0780000016093254, 
    0.034000001847744, 0.0610000006854534, 0.0719999969005585, 
    0.0270000007003546, 0.0850000008940697, 0.0599999986588955, 
    0.0370000004768372, 0.0549999997019768, 0.0790000036358833, 
    0.128000006079674, 0.0439999997615814, 0.0309999994933605, 
    0.0359999984502792, 0.00800000037997961, 0.00300000002607703, 
    0.00800000037997961 ;

 aerosol_optical_depth_8_ = 0.0109999999403954, 0.0270000007003546, 
    0.017000000923872, 0.0430000014603138, 0.025000000372529, 
    0.00899999961256981, 0.0280000008642673, 0.0299999993294477, 
    0.0230000000447035, 0.0309999994933605, 0.0160000007599592, 
    0.0489999987185001, 0.0160000007599592, 0.0230000000447035, 
    0.00899999961256981, 0.0719999969005585, 0.028999999165535, 
    0.0160000007599592, 0.0179999992251396, 0.00400000018998981, 
    0.0130000002682209, 0.0570000000298023, 0.0260000005364418, 
    0.0020000000949949, 0.0230000000447035, 0.00800000037997961, 
    0.00600000005215406, 0.00400000018998981, 0.00300000002607703, 
    0.00100000004749745, 0.00300000002607703, 0.0020000000949949, 
    0.00800000037997961, 0.0230000000447035, 0.0439999997615814, 
    0.0209999997168779, 0.0219999998807907, 0.0769999995827675, 
    0.0140000004321337, 0.0219999998807907, 0.0219999998807907, 
    0.00700000021606684, 0.00899999961256981, 0.00999999977648258, 
    0.0450000017881393, 0.0390000008046627, 0.0350000001490116, 
    0.028999999165535, 0.00300000002607703, 0.00700000021606684, 
    0.00400000018998981, 0.025000000372529, 0.00800000037997961, 
    0.00800000037997961, 0.00700000021606684, 0.0189999993890524, 
    0.00800000037997961, 0.0120000001043081, 0.00800000037997961, 
    0.00800000037997961, 0.0130000002682209, 0.0509999990463257, 
    0.0189999993890524, 0.0020000000949949, 0.00999999977648258, 
    0.0280000008642673, 0, 0.017000000923872, 0.0189999993890524, 
    0.00400000018998981, 0.00600000005215406, 0.00800000037997961, 
    0.0199999995529652, 0.0120000001043081, 0.0120000001043081, 
    0.0140000004321337, 0.00899999961256981, 0.0529999993741512, 
    0.0130000002682209, 0.0149999996647239, 0.0970000028610229, 
    0.00800000037997961, 0.0299999993294477, 0.0710000023245811, 
    0.0209999997168779, 0.0320000015199184, 0.0379999987781048, 
    0.017000000923872, 0.0509999990463257, 0.0370000004768372, 
    0.0199999995529652, 0.034000001847744, 0.0719999969005585, 
    0.0659999996423721, 0.0230000000447035, 0.0270000007003546, 
    0.0320000015199184, 0.00499999988824129, 0.0020000000949949, 
    0.00700000021606684 ;

 aerosol_optical_depth_9_ = 0.00999999977648258, 0.0260000005364418, 
    0.0149999996647239, 0.0419999994337559, 0.0240000002086163, 
    0.00800000037997961, 0.0280000008642673, 0.028999999165535, 
    0.0199999995529652, 0.0299999993294477, 0.0149999996647239, 
    0.0480000004172325, 0.0140000004321337, 0.0199999995529652, 
    0.00800000037997961, 0.0710000023245811, 0.0280000008642673, 
    0.0130000002682209, 0.0149999996647239, 0.00400000018998981, 
    0.0130000002682209, 0.0520000010728836, 0.0209999997168779, 
    0.0020000000949949, 0.0219999998807907, 0.00800000037997961, 
    0.00499999988824129, 0.00400000018998981, 0.00300000002607703, 
    0.00100000004749745, 0.0020000000949949, 0.0020000000949949, 
    0.00800000037997961, 0.0219999998807907, 0.0430000014603138, 
    0.0199999995529652, 0.0209999997168779, 0.0759999975562096, 
    0.0140000004321337, 0.0209999997168779, 0.0209999997168779, 
    0.00700000021606684, 0.00700000021606684, 0.00999999977648258, 
    0.0450000017881393, 0.0379999987781048, 0.0350000001490116, 
    0.0270000007003546, 0.0020000000949949, 0.00600000005215406, 
    0.00400000018998981, 0.0240000002086163, 0.00700000021606684, 
    0.00700000021606684, 0.00600000005215406, 0.0179999992251396, 
    0.00700000021606684, 0.0109999999403954, 0.00700000021606684, 
    0.00700000021606684, 0.0130000002682209, 0.0500000007450581, 
    0.0189999993890524, 0.0020000000949949, 0.00899999961256981, 
    0.0270000007003546, 0, 0.0160000007599592, 0.0179999992251396, 
    0.00400000018998981, 0.00499999988824129, 0.00700000021606684, 
    0.0179999992251396, 0.0109999999403954, 0.0109999999403954, 
    0.0130000002682209, 0.00800000037997961, 0.0520000010728836, 
    0.0130000002682209, 0.0140000004321337, 0.0949999988079071, 
    0.00700000021606684, 0.0270000007003546, 0.0700000002980232, 
    0.0189999993890524, 0.028999999165535, 0.0329999998211861, 
    0.0160000007599592, 0.0469999983906746, 0.034000001847744, 
    0.0179999992251396, 0.0309999994933605, 0.0710000023245811, 
    0.0570000000298023, 0.0179999992251396, 0.0270000007003546, 
    0.0320000015199184, 0.00499999988824129, 0.0020000000949949, 
    0.00700000021606684 ;

 aerosol_optical_depth_10_ = 0.00899999961256981, 0.0260000005364418, 
    0.0130000002682209, 0.0410000011324883, 0.0240000002086163, 
    0.00700000021606684, 0.0270000007003546, 0.0280000008642673, 
    0.017000000923872, 0.028999999165535, 0.0149999996647239, 
    0.0469999983906746, 0.0120000001043081, 0.017000000923872, 
    0.00600000005215406, 0.0700000002980232, 0.0280000008642673, 
    0.0109999999403954, 0.0120000001043081, 0.00300000002607703, 
    0.0130000002682209, 0.046000000089407, 0.017000000923872, 
    0.00100000004749745, 0.0219999998807907, 0.00700000021606684, 
    0.00400000018998981, 0.00400000018998981, 0.0020000000949949, 
    0.00100000004749745, 0.0020000000949949, 0.00100000004749745, 
    0.00700000021606684, 0.0209999997168779, 0.0419999994337559, 
    0.0199999995529652, 0.0209999997168779, 0.0750000029802322, 
    0.0140000004321337, 0.0209999997168779, 0.0209999997168779, 
    0.00600000005215406, 0.00600000005215406, 0.00899999961256981, 
    0.0439999997615814, 0.0370000004768372, 0.034000001847744, 
    0.0230000000447035, 0.0020000000949949, 0.00400000018998981, 
    0.00400000018998981, 0.0230000000447035, 0.00700000021606684, 
    0.00600000005215406, 0.00499999988824129, 0.0179999992251396, 
    0.00600000005215406, 0.0109999999403954, 0.00600000005215406, 
    0.00600000005215406, 0.0120000001043081, 0.0489999987185001, 
    0.0179999992251396, 0.0020000000949949, 0.00899999961256981, 
    0.0260000005364418, 0, 0.0149999996647239, 0.017000000923872, 
    0.00300000002607703, 0.00400000018998981, 0.00600000005215406, 
    0.0160000007599592, 0.00999999977648258, 0.00899999961256981, 
    0.0120000001043081, 0.00600000005215406, 0.0500000007450581, 
    0.0130000002682209, 0.0130000002682209, 0.0930000022053719, 
    0.00700000021606684, 0.0219999998807907, 0.0689999982714653, 
    0.017000000923872, 0.0240000002086163, 0.0280000008642673, 
    0.0140000004321337, 0.0410000011324883, 0.0299999993294477, 
    0.0149999996647239, 0.0270000007003546, 0.0700000002980232, 
    0.0469999983906746, 0.0130000002682209, 0.0260000005364418, 
    0.0309999994933605, 0.00499999988824129, 0.00100000004749745, 
    0.00700000021606684 ;

 aerosol_optical_depth_11_ = 0.00700000021606684, 0.0240000002086163, 
    0.00999999977648258, 0.0390000008046627, 0.0219999998807907, 
    0.00600000005215406, 0.025000000372529, 0.0270000007003546, 
    0.0140000004321337, 0.0280000008642673, 0.0140000004321337, 
    0.0450000017881393, 0.00999999977648258, 0.0140000004321337, 
    0.00300000002607703, 0.0670000016689301, 0.0260000005364418, 
    0.00700000021606684, 0.00700000021606684, 0.0020000000949949, 
    0.0109999999403954, 0.0320000015199184, 0.00999999977648258, 0, 
    0.0189999993890524, 0.00600000005215406, 0.0020000000949949, 
    0.00300000002607703, 0.0020000000949949, 0, 0.00100000004749745, 0, 
    0.00600000005215406, 0.0199999995529652, 0.0399999991059303, 
    0.0179999992251396, 0.0189999993890524, 0.0719999969005585, 
    0.0130000002682209, 0.0189999993890524, 0.0189999993890524, 
    0.00499999988824129, 0.00400000018998981, 0.00899999961256981, 
    0.0419999994337559, 0.0350000001490116, 0.0320000015199184, 
    0.0160000007599592, 0, 0.0020000000949949, 0.00300000002607703, 
    0.0199999995529652, 0.00700000021606684, 0.00499999988824129, 
    0.00300000002607703, 0.017000000923872, 0.00499999988824129, 
    0.00999999977648258, 0.00499999988824129, 0.00400000018998981, 
    0.0109999999403954, 0.0469999983906746, 0.017000000923872, 
    0.0020000000949949, 0.00700000021606684, 0.0230000000447035, 0, 
    0.0130000002682209, 0.0130000002682209, 0.00300000002607703, 
    0.00300000002607703, 0.00400000018998981, 0.0109999999403954, 
    0.00800000037997961, 0.00499999988824129, 0.00999999977648258, 
    0.00400000018998981, 0.0430000014603138, 0.0109999999403954, 
    0.00999999977648258, 0.0820000022649765, 0.00499999988824129, 
    0.0140000004321337, 0.0659999996423721, 0.0149999996647239, 
    0.0189999993890524, 0.0209999997168779, 0.0120000001043081, 
    0.0350000001490116, 0.025000000372529, 0.0120000001043081, 
    0.0230000000447035, 0.0670000016689301, 0.0350000001490116, 
    0.00499999988824129, 0.0240000002086163, 0.028999999165535, 
    0.00400000018998981, 0.00100000004749745, 0.00600000005215406 ;

 aerosol_optical_depth_err_1_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_2_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_3_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_4_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 0, 
    25.6410255432129, 0, 25.6410255432129, 0, 0, 0, 0, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 0, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 0, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 0, 25.6410255432129, 0, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 25.6410255432129, 0, 
    25.6410255432129, 25.6410255432129, 0, 15.151515007019, 15.151515007019, 
    0, 25.6410255432129, 25.6410255432129, 0, 25.6410255432129, 
    25.6410255432129, 0, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 0, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 8.5470085144043, 
    15.151515007019, 8.5470085144043, 8.5470085144043, 15.151515007019, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 25.6410255432129, 15.151515007019, 
    15.151515007019, 0, 0, 0 ;

 aerosol_optical_depth_err_5_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_6_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_7_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_8_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_9_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_10_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_err_11_ = 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 8.5470085144043, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    15.151515007019, 15.151515007019, 15.151515007019, 8.5470085144043, 
    15.151515007019, 15.151515007019, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 15.151515007019, 25.6410255432129, 
    25.6410255432129, 15.151515007019, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019, 25.6410255432129, 25.6410255432129, 
    15.151515007019, 25.6410255432129, 25.6410255432129, 15.151515007019, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 25.6410255432129, 25.6410255432129, 25.6410255432129, 
    25.6410255432129, 8.5470085144043, 15.151515007019, 8.5470085144043, 
    8.5470085144043, 15.151515007019, 8.5470085144043, 8.5470085144043, 
    8.5470085144043, 8.5470085144043, 8.5470085144043, 8.5470085144043, 
    25.6410255432129, 15.151515007019, 15.151515007019, 15.151515007019, 
    15.151515007019, 15.151515007019 ;

 aerosol_optical_depth_qc_1_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_2_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_3_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_4_ = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 
    1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1 ;

 aerosol_optical_depth_qc_5_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_6_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_7_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_8_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_9_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_10_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 aerosol_optical_depth_qc_11_ = -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, 
    -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0, -0 ;

 obs_minus_forecast_unadjusted_1_ = -0.0451268665492535, -0.0514005646109581, 
    0.0123418401926756, -0.0150858573615551, -0.000782416725996882, 
    0.0204685106873512, -0.00418132217600942, 0.0023959104437381, 
    0.1315878033638, 0.023490784689784, -0.00817140284925699, 
    0.054369255900383, 0.0918733179569244, 0.139873817563057, 
    0.0364200249314308, 0.0994362086057663, 0.0338680930435658, 
    0.056239414960146, 0.0539132691919804, 0.0327430106699467, 
    0.00984406471252441, 0.127236023545265, 0.104852594435215, 
    0.0304616000503302, 0.0505893267691135, 0.00516735669225454, 
    0.0192893147468567, 0.0124927368015051, 0.0396594852209091, 
    0.0141699584200978, 0.0306340269744396, 0.0337680950760841, 
    0.0220068302005529, -0.00145220872946084, 0.0530058443546295, 
    0.0210065227001905, 0.0211105849593878, 0.110443413257599, 
    -0.0181664619594812, 0.00203269999474287, 0.0251768119633198, 
    0.0576558150351048, 0.0271848421543837, -0.00542710768058896, 
    0.0409991852939129, 0.0519946776330471, 0.0413541533052921, 
    0.0882418751716614, 0.0509200766682625, 0.0349812544882298, 
    -0.0132404593750834, 0.0279405787587166, -0.00626907683908939, 
    0.0198537409305573, 0.0303867068141699, 0.0184622164815664, 
    0.0639379471540451, 0.00685370899736881, 0.0703121423721313, 
    0.0604482777416706, 0.00212568929418921, 0.00267945160157979, 
    -0.0110704842954874, -0.0255769342184067, 0.0536772198975086, 
    0.102774254977703, -0.01972253061831, 0.0529498867690563, 
    0.00765555119141936, -0.00586831988766789, 0.059288777410984, 
    0.0754664242267609, 0.054257158190012, 0.0250366721302271, 
    0.0254146754741669, 0.0198678690940142, 0.0296585224568844, 
    0.0460681989789009, -0.0227178242057562, 0.110819108784199, 
    0.28352677822113, 0.0681991949677467, 0.215123578906059, 
    0.0904238522052765, 0.0984112173318863, 0.207311049103737, 
    0.235537514090538, 0.0722658708691597, 0.292766630649567, 
    0.188326880335808, 0.100323088467121, 0.163437142968178, 
    0.0802522972226143, 0.423990517854691, 0.0795848667621613, 
    0.0172024555504322, 0.0180104412138462, 0.0088355727493763, 
    -0.0127789843827486, -0.0114837111905217 ;

 obs_minus_forecast_unadjusted_2_ = -0.0514699555933475, -0.0518817566335201, 
    0.00204957369714975, -0.0165077894926071, -0.000567531737033278, 
    0.0155584653839469, -0.00478859432041645, 0.00155591277871281, 
    0.11651649326086, 0.0224743410944939, -0.00818257033824921, 
    0.0511443242430687, 0.0814196467399597, 0.123446978628635, 
    0.0322723016142845, 0.0951621159911156, 0.0324306562542915, 
    0.0501748770475388, 0.0487993061542511, 0.0252879057079554, 
    0.00745825888589025, 0.114743143320084, 0.0973611399531364, 
    0.0228949338197708, 0.0430278219282627, 0.00252776080742478, 
    0.0165981091558933, 0.00882535800337791, 0.0318808630108833, 
    0.0113220224156976, 0.0247906967997551, 0.0278704911470413, 
    0.0180985946208239, -0.00140354689210653, 0.0506662391126156, 
    0.0206190142780542, 0.0197775326669216, 0.104939669370651, 
    -0.0188014172017574, 0.000306015455862507, 0.0245261285454035, 
    0.0482115782797337, 0.023810900747776, -0.00564074888825417, 
    0.0389619655907154, 0.0494706258177757, 0.0386412441730499, 
    0.0776419639587402, 0.0414761826395988, 0.0305857844650745, 
    -0.0134533550590277, 0.0252382513135672, -0.00690770614892244, 
    0.0173214115202427, 0.0268932972103357, 0.0178143195807934, 
    0.0532990545034409, 0.00646654842421412, 0.0586433261632919, 
    0.0518133379518986, 0.00188912183512002, -0.00080350146163255, 
    -0.0120203578844666, -0.0251881554722786, 0.0449930429458618, 
    0.0891826078295708, -0.0191330946981907, 0.0438163988292217, 
    0.0076404963620007, -0.00850840099155903, 0.0486026406288147, 
    0.0628572925925255, 0.0477540716528893, 0.0227341931313276, 
    0.0238059610128403, 0.0182700455188751, 0.0251532252877951, 
    0.0447224341332912, -0.0230644233524799, 0.0938787907361984, 
    0.251612424850464, 0.0572254434227943, 0.185250476002693, 
    0.0860750377178192, 0.0860761776566505, 0.183913201093674, 
    0.209376573562622, 0.062092624604702, 0.259289979934692, 
    0.164054319262505, 0.0862610563635826, 0.142427667975426, 
    0.0763518586754799, 0.379154592752457, 0.0751056000590324, 
    0.0161906033754349, 0.016968309879303, 0.00633796071633697, 
    -0.0133090689778328, -0.0108024505898356 ;

 obs_minus_forecast_unadjusted_3_ = -0.0572427920997143, -0.0528510361909866, 
    -0.00968863628804684, -0.0194240566343069, -0.00201546214520931, 
    0.00993345957249403, -0.00602543540298939, 3.40369588229805e-05, 
    0.0976773872971535, 0.0197211317718029, -0.00891093257814646, 
    0.0471259951591492, 0.0681001842021942, 0.105168960988522, 
    0.0263474602252245, 0.0880808606743813, 0.0291454903781414, 
    0.0423659607768059, 0.0429346039891243, 0.0169736985117197, 
    0.00423255609348416, 0.101382061839104, 0.0869989916682243, 
    0.0144512327387929, 0.0345895811915398, -0.00200591469183564, 
    0.0129982074722648, 0.00425512017682195, 0.0241675078868866, 
    0.00751860439777374, 0.0189915634691715, 0.0210040938109159, 
    0.014220068231225, -0.00304800015874207, 0.0465362817049026, 
    0.0183910857886076, 0.0186217110604048, 0.0975835025310516, 
    -0.0202432498335838, -0.00126866856589913, 0.0219798851758242, 
    0.0379101745784283, 0.0206001028418541, -0.00564092118293047, 
    0.0352240763604641, 0.0450815036892891, 0.0350408293306828, 
    0.0651676803827286, 0.0311770476400852, 0.0263450015336275, 
    -0.0124665573239326, 0.0216651782393456, -0.00741745578125119, 
    0.014904017560184, 0.0235186535865068, 0.0152804534882307, 
    0.042754091322422, 0.00622690469026566, 0.0470636785030365, 
    0.0412702672183514, 0.000872796576004475, -0.00590083887800574, 
    -0.0125996097922325, -0.0246519204229116, 0.035415206104517, 
    0.0746960490942001, -0.019372059032321, 0.0339277163147926, 
    0.00690369121730328, -0.0100114429369569, 0.0370156206190586, 
    0.0503543801605701, 0.0393957309424877, 0.0196242518723011, 
    0.0223024655133486, 0.0157848112285137, 0.0208065789192915, 
    0.0425744764506817, -0.0222050156444311, 0.075963631272316, 
    0.216728821396828, 0.0452718175947666, 0.152418568730354, 
    0.078958585858345, 0.071940504014492, 0.156697243452072, 
    0.177492320537567, 0.0501766316592693, 0.22098246216774, 
    0.137045413255692, 0.0705393403768539, 0.117758892476559, 
    0.0697754546999931, 0.325650066137314, 0.0687920749187469, 
    0.0144503358751535, 0.0142309591174126, 0.00299508054740727, 
    -0.0136864418163896, -0.0109173059463501 ;

 obs_minus_forecast_unadjusted_4_ = -0.0876630246639252, -0.0766100659966469, 
    -0.0137223722413182, -0.0161074865609407, -0.0266869068145752, 
    -0.0180435683578253, -0.0304070170968771, -0.0247520990669727, 
    0.0959437415003777, -0.00543440552428365, -0.0319890417158604, 
    0.0509844832122326, 0.0602274127304554, 0.102386832237244, 
    -0.00206604576669633, 0.102859370410442, 0.0042049209587276, 
    0.0111459568142891, 0.0126394331455231, -0.0130094168707728, 
    -0.0206204820424318, 0.0653293877840042, 0.0519383512437344, 
    -0.0157071501016617, 0.00343771907500923, -0.02429274097085, 
    -0.0123920012265444, -0.017091266810894, -0.00639648921787739, 
    -0.0081823356449604, -0.00770540256053209, -0.00878919940441847, 
    -0.00958963017910719, -0.0269803404808044, 0.0473397858440876, 
    -0.00647699553519487, -0.00613486021757126, 0.113507255911827, 
    -0.0432279594242573, -0.0264837834984064, -0.00332851381972432, 
    0.00393130350857973, -0.00624256860464811, -0.0211606100201607, 
    0.0374634228646755, 0.0435203462839127, 0.0325418002903461, 
    0.0309796277433634, -0.00179491424933076, -0.00154701550491154, 
    -0.018028948456049, -0.00460263201966882, -0.0196324530988932, 
    -0.0102531677111983, -0.00358675280585885, -0.00899145286530256, 
    0.00842281896620989, -0.0126794194802642, 0.0116859385743737, 
    0.00793467927724123, -0.0196521822363138, -0.00045362624223344, 
    -0.0363354384899139, -0.027768274769187, 0.00208305194973946, 
    0.0364484339952469, -0.0182199999690056, 0.00159288675058633, 
    -0.0162030942738056, -0.0251908227801323, 0.00265602744184434, 
    0.0130947744473815, 0.00936655327677727, -0.00704987626522779, 
    -0.00196063867770135, -0.00844165962189436, -0.00717234006151557, 
    0.0178874414414167, -0.0358635410666466, 0.0351077057421207, 
    0.156917676329613, 0.0103679765015841, 0.0946840718388557, 
    0.0929426401853561, 0.0643331557512283, 0.16353203356266, 
    0.158235639333725, 0.042457289993763, 0.195053562521935, 
    0.141334176063538, 0.0681301057338715, 0.120521560311317, 
    0.0839342698454857, 0.278896242380142, 0.0378556586802006, 
    -0.0106741804629564, -0.0108178136870265, -0.0179947055876255, 
    -0.0197149161249399, -0.0215715728700161 ;

 obs_minus_forecast_unadjusted_5_ = -0.0708276778459549, -0.0524899512529373, 
    -0.0375378504395485, -0.0231127608567476, -0.00367669016122818, 
    -0.00265276455320418, -0.00792767014354467, -0.00389652349986136, 
    0.0481566078960896, 0.0146799013018608, -0.00865704938769341, 
    0.0360907092690468, 0.0347157567739487, 0.0539995208382607, 
    0.0105826510116458, 0.071729376912117, 0.0229984875768423, 
    0.0201697610318661, 0.0225754044950008, -0.000280729407677427, 
    -0.00166592409368604, 0.0709302723407745, 0.054511483758688, 
    -0.00425602030009031, 0.0148963816463947, -0.00901100318878889, 
    0.00366972456686199, -0.00495809502899647, 0.00537237757816911, 
    -0.000654340838082135, 0.00482406280934811, 0.00458861794322729, 
    0.0047639892436564, -0.00434295041486621, 0.0362733639776707, 
    0.0144189978018403, 0.0149569800123572, 0.0782887935638428, 
    -0.0219909753650427, -0.00670956587418914, 0.016904329881072, 
    0.01363789383322, 0.00970324221998453, -0.00462430808693171, 
    0.0266438722610474, 0.0355780720710754, 0.0260131787508726, 
    0.0384488999843597, 0.00793613772839308, 0.0123099023476243, 
    -0.0106248538941145, 0.0119057381525636, -0.00813706032931805, 
    0.00814877543598413, 0.0118748620152473, 0.0113347871229053, 
    0.0175469685345888, 0.00511796912178397, 0.0187381561845541, 
    0.0180402547121048, 0.000888232025317848, -0.0148733928799629, 
    -0.0131483534350991, -0.0230246912688017, 0.0123081691563129, 
    0.0407087355852127, -0.0162044614553452, 0.0134603856131434, 
    0.00507281767204404, -0.014573585242033, 0.0108274705708027, 
    0.018360773101449, 0.0220632683485746, 0.0102121671661735, 
    0.0162890776991844, 0.00989237986505032, 0.00670227687805891, 
    0.0372259542346001, -0.0194118749350309, 0.0343980267643929, 
    0.135279566049576, 0.0165955070406199, 0.0751764923334122, 
    0.0629765391349792, 0.0345516130328178, 0.0829820483922958, 
    0.091376967728138, 0.0217655170708895, 0.1199636682868, 
    0.0675864666700363, 0.0293741375207901, 0.0566677041351795, 
    0.0557612888514996, 0.17482428252697, 0.0447868071496487, 
    0.010561971925199, 0.00970939919352531, -0.00318795838393271, 
    -0.0139314020052552, -0.0091950511559844 ;

 obs_minus_forecast_unadjusted_6_ = -0.0726091042160988, -0.0507462844252586, 
    -0.0425966344773769, -0.022505609318614, -0.003422393463552, 
    -0.00479604722931981, -0.0084111150354147, -0.0036960793659091, 
    0.0366703718900681, 0.014394081197679, -0.00877293758094311, 
    0.0345044247806072, 0.0265973135828972, 0.0419682152569294, 
    0.00702539412304759, 0.0679899528622627, 0.0219872761517763, 
    0.0148507570847869, 0.0172141790390015, -0.00331078027375042, 
    -0.00257105776108801, 0.0648211464285851, 0.0453784242272377, 
    -0.00743406265974045, 0.011717801913619, -0.0102619733661413, 
    0.0012742878170684, -0.00631593354046345, 0.00181333487853408, 
    -0.00235157646238804, 0.00212510023266077, 0.00181186851114035, 
    0.0029776229057461, -0.00425708666443825, 0.0346407406032085, 
    0.0144501021131873, 0.0140973972156644, 0.0752697885036469, 
    -0.0214752033352852, -0.00648812158033252, 0.0156160360202193, 
    0.00856489967554808, 0.006764923222363, -0.00421703280881047, 
    0.0256502162665129, 0.0344618484377861, 0.0248403251171112, 
    0.0323054865002632, 0.00388298486359417, 0.00832062587141991, 
    -0.00931940693408251, 0.00988166127353907, -0.00722676469013095, 
    0.00590889807790518, 0.00965425465255976, 0.0101134842261672, 
    0.0121633494272828, 0.00507805403321981, 0.013319474644959, 
    0.0136389974504709, 0.00029827150865458, -0.0149101316928864, 
    -0.0116776004433632, -0.021929893642664, 0.00903153419494629, 
    0.0343962013721466, -0.0150672225281596, 0.0100541422143579, 
    0.0049058748409152, -0.0155575051903725, 0.00651933718472719, 
    0.0130670154467225, 0.0190217364579439, 0.00845813844352961, 
    0.0139817567542195, 0.00864325929433107, 0.00281618838198483, 
    0.0355794243514538, -0.0179599672555923, 0.0255820974707603, 
    0.119501888751984, 0.0107542397454381, 0.0594718344509602, 
    0.0605230331420898, 0.0268437955528498, 0.0661570131778717, 
    0.0711847767233849, 0.0164165124297142, 0.0970516726374626, 
    0.0533288568258286, 0.0205914471298456, 0.0438653379678726, 
    0.0529519207775593, 0.138050213456154, 0.0379137024283409, 
    0.0103711253032088, 0.00975585170090199, -0.00514479866251349, 
    -0.013879562728107, -0.00884284731000662 ;

 obs_minus_forecast_unadjusted_7_ = -0.0721308439970016, -0.0480394996702671, 
    -0.0456763990223408, -0.0200961846858263, -0.00320959673263133, 
    -0.00621999008581042, -0.00682056834921241, -0.0035085731651634, 
    0.0247527714818716, 0.0147834904491901, -0.00709300069138408, 
    0.0325274392962456, 0.0188068859279156, 0.030310770496726, 
    0.00302942679263651, 0.0647420659661293, 0.0203679222613573, 
    0.00920560397207737, 0.0115351369604468, -0.00692904088646173, 
    -0.00201093452051282, 0.0580807365477085, 0.0345918051898479, 
    -0.01025456096977, 0.00889908988028765, -0.0111431609839201, 
    -0.00185057998169214, -0.00738795101642609, -0.00154209567699581, 
    -0.00390916550531983, -0.000437881040852517, -0.00185108126606792, 
    0.00130405696108937, -0.00325308251194656, 0.0335999615490437, 
    0.0138745559379458, 0.0136779574677348, 0.0706721544265747, 
    -0.0209981594234705, -0.006469642277807, 0.0146490624174476, 
    0.00483932951465249, 0.00423112185671926, -0.00324287475086749, 
    0.0245618745684624, 0.0317074693739414, 0.023127855733037, 
    0.0275582745671272, 0.000192003295524046, 0.00471512321382761, 
    -0.00752271572127938, 0.00842780526727438, -0.00684748496860266, 
    0.00395464804023504, 0.00671036029234529, 0.0102603249251842, 
    0.00801912322640419, 0.00437996536493301, 0.00812952686101198, 
    0.00846333988010883, 0.00126585457473993, -0.0139815434813499, 
    -0.0100512411445379, -0.0202224515378475, 0.00510015152394772, 
    0.0283496119081974, -0.0134444357827306, 0.00728755863383412, 
    0.00449252594262362, -0.014977945946157, 0.00154701294377446, 
    0.00706646731123328, 0.015390869230032, 0.00619290489703417, 
    0.0119512481614947, 0.00770974764600396, -0.000520104949828237, 
    0.0345585830509663, -0.0157945714890957, 0.0168737545609474, 
    0.104844480752945, 0.00502029061317444, 0.0439179427921772, 
    0.0577947869896889, 0.0196736808866262, 0.0488117188215256, 
    0.0507834143936634, 0.0107550164684653, 0.0736015141010284, 
    0.0378803908824921, 0.0118149928748608, 0.0310262888669968, 
    0.0511159524321556, 0.100248135626316, 0.0285635944455862, 
    0.010927869938314, 0.00973719451576471, -0.00563156045973301, 
    -0.0123250838369131, -0.00790724344551563 ;

 obs_minus_forecast_unadjusted_8_ = -0.0618702881038189, -0.035136915743351, 
    -0.0426687598228455, -0.0105187864974141, 0.0016978126950562, 
    -0.00618165358901024, -0.00189255480654538, 0.00164267094805837, 
    0.0105725796893239, 0.0164161343127489, -0.0025224625132978, 
    0.032599613070488, 0.00861128605902195, 0.0144556788727641, 
    -0.00229172594845295, 0.0618747062981129, 0.0206354632973671, 
    0.00182476127520204, 0.00315570598468184, -0.00846936833113432, 
    -0.000118298739835154, 0.0461752526462078, 0.0165206454694271, 
    -0.0132480002939701, 0.00790378078818321, -0.0101512633264065, 
    -0.00559307029470801, -0.00800406001508236, -0.00487275095656514, 
    -0.00474682822823524, -0.00230770907364786, -0.00491465302184224, 
    0.000234066363191232, 0.00131186086218804, 0.0333992056548595, 
    0.0141650978475809, 0.0143376821652055, 0.0671321600675583, 
    -0.0153934210538864, -0.00315304822288454, 0.0142846051603556, 
    0.000767026038374752, 0.00162762345280498, -0.00052885920740664, 
    0.0269317887723446, 0.0307173188775778, 0.0218156110495329, 
    0.0197865478694439, -0.00376367708668113, -5.82309330638964e-05, 
    -0.00438732886686921, 0.00796705670654774, -0.00407625362277031, 
    0.0023799785412848, 0.0020851269364357, 0.0102433385327458, 
    0.00303022703155875, 0.00629594875499606, 0.00304747256450355, 
    0.00336694205179811, 0.0038550766184926, -0.00461427634581923, 
    -0.0037625739350915, -0.0163392927497625, 0.00187392835505307, 
    0.0225766524672508, -0.0094562629237771, 0.00655944878235459, 
    0.00572034856304526, -0.0124669438228011, -0.00272440258413553, 
    0.00149855914060026, 0.0117701040580869, 0.00423803646117449, 
    0.00626386143267155, 0.00731761194765568, -0.00406928872689605, 
    0.0336440242826939, -0.0110246008262038, 0.00774096325039864, 
    0.0898140221834183, -0.00112743722274899, 0.0221334025263786, 
    0.0566084943711758, 0.0110539263114333, 0.0237336903810501, 
    0.0231702551245689, 0.00630902592092752, 0.0433311760425568, 
    0.0213474575430155, 0.0028579467907548, 0.0177678558975458, 
    0.0521081835031509, 0.046242032200098, 0.011825131252408, 
    0.0131290107965469, 0.0133202215656638, -0.00478369882330298, 
    -0.00923401582986116, -0.00412403466179967 ;

 obs_minus_forecast_unadjusted_9_ = -0.0573872849345207, -0.0314043201506138, 
    -0.0400281250476837, -0.00730262883007526, 0.00281065725721419, 
    -0.00564520573243499, 0.000536263221874833, 0.00291766389273107, 
    0.00878699962049723, 0.0168542470782995, -0.00178195489570498, 
    0.0329898931086063, 0.00732117239385843, 0.0122574232518673, 
    -0.00210258550941944, 0.0619331449270248, 0.020475871860981, 
    0.000279332016361877, 0.00162958260625601, -0.00751379551365972, 
    0.00094969553174451, 0.0420151986181736, 0.0123021081089973, 
    -0.0123833725228906, 0.00776672549545765, -0.0092629985883832, 
    -0.00593405542895198, -0.00731134414672852, -0.00439162971451879, 
    -0.00440266635268927, -0.00297863711602986, -0.0046184416860342, 
    0.000535375962499529, 0.00236599124036729, 0.0336623787879944, 
    0.0139923030510545, 0.0142610799521208, 0.0670521706342697, 
    -0.0129901524633169, -0.00212760758586228, 0.0140117835253477, 
    0.0014972286298871, 0.000482673931401223, 0.000697196053806692, 
    0.0289459582418203, 0.0305053070187569, 0.0229304488748312, 
    0.0186819229274988, -0.00399493100121617, -0.000245136849116534, 
    -0.00335011957213283, 0.00836198031902313, -0.00397692481055856, 
    0.00199480797164142, 0.00166830723173916, 0.0100767528638244, 
    0.00254528550431132, 0.00600606389343739, 0.00254211109131575, 
    0.0028474482242018, 0.00500657362863421, -0.000715959758963436, 
    -0.00121953908819705, -0.0148603776469827, 0.00164410809520632, 
    0.0221448596566916, -0.00839197542518377, 0.00690244417637587, 
    0.00634475192055106, -0.011104341596365, -0.00294319749809802, 
    0.0011452678591013, 0.0106771932914853, 0.00425474159419537, 
    0.00586237292736769, 0.00700754625722766, -0.00379149592481554, 
    0.0340643748641014, -0.00935945753008127, 0.00702687026932836, 
    0.0881182923913002, -0.00183147424831986, 0.0194997061043978, 
    0.0571878701448441, 0.0101795857772231, 0.0217280853539705, 
    0.0198408309370279, 0.00671683438122272, 0.040288507938385, 
    0.0200845971703529, 0.002980433171615, 0.0167801566421986, 
    0.0533007495105267, 0.0394205562770367, 0.00801228452473879, 
    0.014762993901968, 0.0153963649645448, -0.0037253494374454, 
    -0.00807503517717123, -0.00284899258986115 ;

 obs_minus_forecast_unadjusted_10_ = -0.0504122376441956, 
    -0.0245508085936308, -0.0353957675397396, -0.00228601391427219, 
    0.00569722894579172, -0.00460773659870028, 0.0028973191510886, 
    0.00511164963245392, 0.00738976150751114, 0.0177633967250586, 
    0.000579369487240911, 0.0339238122105598, 0.00626201182603836, 
    0.0103217093273997, -0.00252558127976954, 0.0623427517712116, 
    0.021596897393465, 0.000229634024435654, 0.000619964150246233, 
    -0.00717237684875727, 0.00243999529629946, 0.0371833145618439, 
    0.00937834847718477, -0.0121263992041349, 0.00901990197598934, 
    -0.00896340329200029, -0.00596779584884644, -0.00629916321486235, 
    -0.00469734892249107, -0.00389553839340806, -0.00249910028651357, 
    -0.00516531569883227, 1.62018056926172e-06, 0.00419320445507765, 
    0.0343699902296066, 0.0150840058922768, 0.0154830487444997, 
    0.0673013404011726, -0.00942134764045477, 0.00090182718122378, 
    0.0150223495438695, 0.00145516917109489, 0.000612210656981915, 
    0.0013505668612197, 0.0307351034134626, 0.0305667165666819, 
    0.0235536377876997, 0.0159282609820366, -0.00297865597531199, 
    -0.00116955942939967, -0.00198122765868902, 0.00940902717411518, 
    -0.00240550166927278, 0.00181115348823369, 0.00142768805380911, 
    0.011240903288126, 0.00223155575804412, 0.00692526903003454, 
    0.00220378744415939, 0.00248269829899073, 0.00551881222054362, 
    0.00558779155835509, 0.00129562756046653, -0.0127016603946686, 
    0.00271610869094729, 0.0219019372016191, -0.00693482859060168, 
    0.00768566271290183, 0.00753572443500161, -0.0101186754181981, 
    -0.00283390516415238, 0.00102884264197201, 0.009923598729074, 
    0.00459327828139067, 0.00466448906809092, 0.00694337207823992, 
    -0.00397674180567265, 0.0340597331523895, -0.00697958515956998, 
    0.00647097872570157, 0.0865774601697922, -0.00136076647322625, 
    0.015039031393826, 0.0583509020507336, 0.00967346597462893, 
    0.0180376470088959, 0.017080994322896, 0.00656759506091475, 
    0.0355578921735287, 0.0184482056647539, 0.00283654732629657, 
    0.015466071665287, 0.055350087583065, 0.0324408039450645, 
    0.00467360485345125, 0.0159816425293684, 0.017269853502512, 
    -0.00225360179319978, -0.00743829971179366, -0.00111067539546639 ;

 obs_minus_forecast_unadjusted_11_ = -0.0343936420977116, 
    -0.0111855128780007, -0.0238563064485788, 0.00885933358222246, 
    0.00948856119066477, -0.00178444001358002, 0.00788496527820826, 
    0.0109446542337537, 0.00738020427525043, 0.0203440710902214, 
    0.00420657498762012, 0.0359831303358078, 0.00603870768100023, 
    0.00933721382170916, -0.00255378964357078, 0.0620158538222313, 
    0.0217350237071514, -9.3420112534659e-06, -0.000479225709568709, 
    -0.00524558825418353, 0.00362401269376278, 0.0257027745246887, 
    0.00465001352131367, -0.00996595434844494, 0.00915791280567646, 
    -0.00669309450313449, -0.00551496911793947, -0.00475148856639862, 
    -0.00303335255011916, -0.00363140483386815, -0.0023338592145592, 
    -0.00492020836099982, 0.000323713989928365, 0.00888668838888407, 
    0.0356665179133415, 0.0151017522439361, 0.0157654080539942, 
    0.0667540803551674, -0.0021825113799423, 0.00598309794440866, 
    0.0151066016405821, 0.00221071345731616, 0.000718844996299595, 
    0.00456967251375318, 0.0344230271875858, 0.0306316930800676, 
    0.0251917224377394, 0.0114990901201963, -0.0030816625803709, 
    -0.00115867715794593, -0.000435693073086441, 0.011064731515944, 
    0.00100152078084648, 0.00235285889357328, 0.000800239620730281, 
    0.0126544134691358, 0.00253297993913293, 0.0075624193996191, 
    0.00247255666181445, 0.00167651812080294, 0.00727727822959423, 
    0.0205733571201563, 0.00741006853058934, -0.00779759651049972, 
    0.00291728950105608, 0.0203403029590845, -0.00404048291966319, 
    0.00899595208466053, 0.00775531213730574, -0.00563188642263412, 
    -0.00144887017086148, 0.000790183374192566, 0.00741982273757458, 
    0.00502113671973348, 0.00219366513192654, 0.00676934514194727, 
    -0.00211016065441072, 0.0314510203897953, -0.00359585322439671, 
    0.00474817585200071, 0.076817013323307, -0.00191353668924421, 
    0.00841706153005362, 0.0596026405692101, 0.0104282544925809, 
    0.0154177928343415, 0.0142997782677412, 0.00789137743413448, 
    0.0318893976509571, 0.0180265679955482, 0.00520467385649681, 
    0.0164368320256472, 0.0586156956851482, 0.0266273282468319, 
    0.000118352159915958, 0.0183297507464886, 0.0210930164903402, 
    -0.000241096131503582, -0.00398682337254286, 0.00130409409757704 ;

 surface_air_pressure_1_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_2_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_3_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_4_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_5_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_6_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_7_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_8_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_9_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_10_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;

 surface_air_pressure_11_ = 980.932556152344, 984.017822265625, 
    984.982543945312, 982.346313476562, 994.665405273438, 994.248107910156, 
    996.576354980469, 990.959777832031, 996.01708984375, 995.175659179688, 
    996.381896972656, 993.692260742188, 1000.41412353516, 997.042724609375, 
    1007.10052490234, 1003.36187744141, 1001.7470703125, 1008.87963867188, 
    1009.05108642578, 1011.49389648438, 1011.0693359375, 1011.79718017578, 
    1011.57501220703, 1014.71417236328, 1014.58947753906, 1011.91833496094, 
    1015.08532714844, 1014.85308837891, 1014.92962646484, 1015.86175537109, 
    1015.46820068359, 1015.83404541016, 1015.77618408203, 995.594177246094, 
    1002.33673095703, 1005.58447265625, 1002.43548583984, 994.52294921875, 
    995.903930664062, 995.399597167969, 1006.64398193359, 1007.84222412109, 
    1005.51977539062, 1003.01422119141, 1001.32177734375, 996.175720214844, 
    1001.88757324219, 1005.04370117188, 1007.20288085938, 1005.59466552734, 
    1004.49029541016, 1006.24487304688, 1006.45104980469, 1007.44946289062, 
    1005.73065185547, 1007.30517578125, 1008.67333984375, 1003.47235107422, 
    1009.26696777344, 1007.47442626953, 1003.81182861328, 1002.2744140625, 
    1001.89489746094, 1007.62396240234, 1009.44439697266, 1008.77801513672, 
    1006.5205078125, 1004.82385253906, 1001.98596191406, 1009.3037109375, 
    1010.21520996094, 1010.3154296875, 1008.36065673828, 1003.72418212891, 
    1011.90881347656, 1011.95220947266, 1011.50756835938, 1011.04241943359, 
    1011.27447509766, 1015.15985107422, 1014.58081054688, 1014.546875, 
    1011.92486572266, 947.990295410156, 943.647766113281, 917.438903808594, 
    915.066833496094, 955.02880859375, 905.614929199219, 910.375061035156, 
    959.581787109375, 960.525756835938, 999.414306640625, 998.867614746094, 
    992.503540039062, 999.0732421875, 999.875305175781, 991.412780761719, 
    997.08984375, 997.532836914062 ;
}
