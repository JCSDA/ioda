netcdf sample_hofx_output_amsua_n19 {
dimensions:
	Channel = 15 ;
	Location = UNLIMITED ; // (17 currently)
variables:
	int Channel(Channel) ;
		Channel:suggested_chunk_dim = 100LL ;
	int Location(Location) ;
		Location:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
data:

 Channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

group: EffectiveError {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5 ;
  } // group EffectiveError

group: GsiFinalObsError {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  -3.368795e+38, -3.368795e+38, -3.368795e+38, -3.368795e+38, 
      -3.368795e+38, -3.368795e+38, 0.2321299, 0.2500168, 0.2500067, 
      0.3500332, 0.4001701, 0.5510925, 0.8075905, 3.136678, -3.368795e+38,
  7.346854, 8.660736, 6.638414, 1.652725, 0.4421597, 0.2319498, 0.2300027, 
      0.2500024, 0.250006, 0.35003, 0.4001538, 0.5509878, 0.8068625, 
      3.123467, 16.91724,
  -3.368795e+38, -3.368795e+38, -3.368795e+38, -3.368795e+38, 
      -3.368795e+38, 0.2311433, 0.2300089, 0.2500034, 0.2500082, 0.3500407, 
      0.4002089, 0.5513419, 0.809324, 3.168164, -3.368795e+38,
  5.185898, 7.67515, 6.818451, 1.567033, 0.7223942, 0.2301599, 0.2300035, 
      -3.368795e+38, 0.2500061, 0.3500302, 0.4001551, 0.5509965, 0.8069223, 
      3.124473, 15.5676,
  -3.368795e+38, -3.368795e+38, -3.368795e+38, -3.368795e+38, 
      -3.368795e+38, 0.2381857, 0.230148, 0.250003, 0.2500059, 0.3500291, 
      0.4001494, 0.5509597, 0.8066677, 3.120001, -3.368795e+38,
  -3.368795e+38, -3.368795e+38, -3.368795e+38, -3.368795e+38, 
      -3.368795e+38, 0.2321259, 0.230022, -3.368795e+38, 0.2500065, 
      0.3500322, 0.4001652, 0.5510617, 0.8073763, 3.132789, -3.368795e+38,
  7.04636, 7.110909, 4.415892, 1.41418, 0.4979441, 0.2354702, 0.2300803, 
      -3.368795e+38, 0.2500058, 0.3500288, 0.4001477, 0.550949, 0.8065947, 
      3.118784, 6.844889,
  7.658558, 8.355218, 7.22888, 1.575394, 0.4435094, 0.2300648, 0.2300024, 
      -3.368795e+38, 0.2500062, 0.3500306, 0.4001569, 0.5510077, 0.8070011, 
      3.126005, 17.5889,
  -3.368795e+38, -3.368795e+38, -3.368795e+38, -3.368795e+38, 
      -3.368795e+38, 0.6543594, 0.2395212, -3.368795e+38, 0.2500066, 
      0.350033, 0.400169, 0.5510858, 0.8075445, 3.135873, -3.368795e+38,
  3.45505, 3.596697, 2.430949, 0.7033065, 0.3388874, 0.2300125, 0.2300027, 
      -3.368795e+38, 0.2500075, 0.3500353, 0.4001774, 0.5511349, 0.80788, 
      3.142086, 4.500139,
  -3.368795e+38, -3.368795e+38, -3.368795e+38, -3.368795e+38, 
      -3.368795e+38, -3.368795e+38, 0.2300046, -3.368795e+38, 0.2500059, 
      0.3500295, 0.4001511, 0.5509709, 0.8067449, 3.121392, -3.368795e+38,
  4.011971, 4.844544, 3.672333, 0.9819183, 0.3468478, 0.2300902, 
      -3.368795e+38, 0.2500024, 0.2500058, 0.3500288, 0.4001475, 0.5509479, 
      0.8065864, 3.118601, 7.93484,
  4.687037, 4.723842, 3.49545, 0.9800412, 0.4253824, 0.2300886, 0.2300027, 
      -3.368795e+38, 0.2500058, 0.3500288, 0.4001476, 0.5509483, 0.8065891, 
      3.11865, 6.206744,
  4.107744, 4.883582, 3.686612, 0.976931, 0.3371014, 0.2300803, 0.230003, 
      -3.368795e+38, 0.2500063, 0.3500296, 0.400149, 0.5509537, 0.806621, 
      3.119228, 8.129551,
  44.45079, 52.53493, 39.16499, 8.894402, 1.291667, 0.2439306, 0.2300024, 
      -3.368795e+38, 0.2500059, 0.3500291, 0.4001494, 0.5509596, 0.806667, 
      3.119985, 61.87202,
  8.41289, 6.911407, 5.486331, 1.309232, 0.4173437, 0.2300978, 0.2300033, 
      0.2500029, 0.2500062, 0.3500291, 0.4001465, 0.5509372, 0.8065058, 
      3.117133, 10.64392,
  -3.368795e+38, -3.368795e+38, -3.368795e+38, -3.368795e+38, 
      -3.368795e+38, 0.2325132, -3.368795e+38, -3.368795e+38, 0.2500056, 
      0.3500277, 0.4001419, 0.5509118, 0.8063363, 3.114146, -3.368795e+38 ;
  } // group GsiFinalObsError

group: GsiHofX {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  176.7687, 174.3334, 195.1922, 214.461, 221.9126, 220.6024, 216.2201, 
      213.0971, 209.6615, 207.6245, 207.8295, 212.1449, 220.7394, 233.5807, 
      181.5459,
  172.2683, 164.0731, 228.8642, 257.6087, 253.9831, 238.99, 226.9764, 
      217.6271, 211.1901, 214.9771, 220.9799, 228.1783, 236.7679, 245.555, 
      234.995,
  288.1978, 288.2496, 282.2845, 269.4221, 254.1952, 234.2566, 220.6119, 
      210.1823, 204.6339, 213.1582, 224.6517, 235.3238, 246.2464, 255.1458, 
      279.0576,
  144.841, 146.998, 213.4474, 246.4555, 245.7055, 234.1104, 225.9846, 
      221.1559, 219.5439, 220.1791, 222.3776, 227.8584, 235.7984, 243.4688, 
      201.5242,
  283.6747, 283.5335, 282.6513, 274.2106, 261.54, 242.507, 227.9962, 
      215.4803, 203.5544, 209.6569, 221.0405, 233.3168, 244.0887, 253.5977, 
      285.5602,
  294.9745, 295.3118, 289.1847, 275.1755, 259.3676, 239.5334, 226.5192, 
      216.3309, 206.6951, 212.7114, 223.2303, 233.0237, 240.919, 248.2065, 
      289.5423,
  257.1417, 254.4036, 254.0532, 252.6951, 244.3344, 231.0919, 222.6275, 
      217.2267, 213.7644, 215.3497, 221.063, 230.0097, 242.2139, 255.3442, 
      249.5818,
  173.791, 162.3867, 229.4941, 261.2972, 256.8979, 240.4063, 227.2521, 
      216.5718, 207.5558, 212.7589, 220.9984, 229.0764, 238.0735, 247.6797, 
      239.072,
  252.897, 251.7748, 252.1441, 251.8353, 245.6719, 232.8181, 222.6957, 
      215.5074, 212.0912, 215.3495, 222.4933, 231.6127, 241.3997, 251.493, 
      247.6844,
  166.2597, 163.1058, 229.3272, 252.6007, 245.6657, 230.9379, 221.262, 
      215.1953, 214.4513, 216.8949, 220.7201, 228.6471, 241.2698, 255.469, 
      221.0255,
  145.6847, 153.3012, 214.5339, 243.2, 243.2445, 234.7629, 228.3755, 
      224.0211, 217.3138, 212.9561, 210.1373, 211.8351, 219.1982, 231.8862, 
      203.4303,
  197.9114, 169.8556, 233.5681, 264.3528, 259.7067, 242.2487, 227.9277, 
      215.7158, 204.2333, 210.3923, 221.8543, 234.4745, 246.2723, 256.235, 
      250.4558,
  189.9944, 165.0524, 230.0302, 263.3905, 259.6016, 242.3235, 227.8974, 
      215.5627, 203.7496, 209.5112, 221.4615, 235.0051, 246.9802, 256.2195, 
      244.8104,
  187.059, 166.8722, 230.8825, 259.2189, 254.1045, 237.9813, 225.8561, 
      216.6842, 210.6434, 215.3035, 224.3548, 234.8271, 245.3712, 255.9125, 
      238.8376,
  181.0434, 183.0752, 242.8816, 256.6268, 251.0137, 237.5273, 227.2836, 
      219.4202, 212.3235, 213.1557, 216.9743, 224.1078, 233.9842, 244.3832, 
      261.1627,
  166.2495, 154.6008, 222.1374, 260.1763, 257.6862, 241.1478, 227.6112, 
      216.7068, 207.3217, 212.2987, 222.0651, 232.5003, 243.2285, 254.5276, 
      223.9976,
  227.3031, 205.3571, 222.5137, 243.7873, 241.6514, 231.5924, 225.0807, 
      221.408, 219.4319, 219.2683, 221.4535, 227.9565, 238.834, 251.822, 
      187.7648 ;
  } // group GsiHofX

group: GsiHofXBc {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  176.5981, 175.5688, 197.1707, 216.2307, 221.8295, 219.6692, 215.2943, 
      212.8763, 208.979, 206.9435, 207.3559, 212.0341, 221.3427, 234.7563, 
      181.2727,
  173.3767, 164.9576, 229.3039, 256.9185, 253.3876, 238.1089, 225.7654, 
      218.3584, 210.5098, 214.4884, 220.5381, 227.9937, 236.9303, 246.0429, 
      235.6887,
  286.7413, 287.1906, 281.3291, 267.8255, 252.3729, 232.8801, 219.1333, 
      212.0711, 203.8756, 212.7783, 224.1915, 235.1262, 246.4018, 255.7163, 
      278.2574,
  146.2813, 148.4597, 214.1299, 245.9193, 245.195, 233.2915, 224.9408, 
      220.4554, 218.8906, 219.5924, 221.923, 227.6917, 235.9309, 244.0675, 
      202.2662,
  283.818, 282.2456, 282.7508, 274.4879, 261.1007, 241.6244, 226.7672, 
      216.315, 202.9272, 209.3798, 220.7717, 233.2777, 244.3311, 254.1851, 
      285.1019,
  293.9211, 293.4003, 288.8949, 274.9675, 258.666, 238.4777, 225.1962, 
      217.5707, 205.8609, 212.2239, 222.7153, 232.6782, 240.7962, 248.5411, 
      289.0827,
  256.986, 254.1251, 254.3117, 252.9867, 243.9593, 230.2301, 221.5174, 
      217.0427, 213.0219, 214.7782, 220.6278, 229.924, 242.6752, 255.7997, 
      248.812,
  174.7889, 163.0416, 230.1367, 260.5786, 256.1994, 239.475, 226.0994, 
      217.6415, 206.9716, 212.4314, 220.6693, 228.993, 238.3879, 248.2577, 
      240.0834,
  252.4661, 252.1985, 253.2206, 253.0155, 245.3248, 231.8046, 221.6635, 
      215.7266, 211.4694, 214.912, 222.1561, 231.5531, 241.7478, 252.0677, 
      247.2725,
  165.7463, 162.8309, 228.654, 251.1478, 244.464, 229.5722, 219.8194, 
      215.5402, 213.3631, 215.8947, 219.8351, 228.1533, 241.4343, 255.5746, 
      222.3541,
  147.2043, 155.2341, 215.7403, 242.9578, 242.8174, 233.959, 227.3614, 
      224.2652, 216.6357, 212.2103, 209.6077, 211.6612, 219.7556, 233.1066, 
      204.3089,
  198.9599, 170.1957, 234.0898, 263.6622, 259.0507, 241.3554, 226.7333, 
      216.6103, 203.6411, 210.1511, 221.6207, 234.5059, 246.604, 256.8594, 
      251.1308,
  190.9139, 165.3457, 230.3424, 262.65, 258.9651, 241.4346, 226.6351, 
      216.4277, 203.0678, 209.2006, 221.183, 234.9776, 247.1872, 256.7917, 
      245.4137,
  187.8503, 167.0183, 231.1406, 258.4549, 253.4742, 237.0778, 224.6344, 
      217.4172, 209.942, 214.872, 223.973, 234.7043, 245.6248, 256.3659, 
      239.4382,
  182.1543, 183.7701, 243.3075, 256.0046, 250.4601, 236.677, 226.1429, 
      220.0346, 211.6548, 212.6052, 216.5654, 224.0205, 234.3372, 244.9175, 
      261.4656,
  167.5791, 155.6027, 222.6802, 259.4971, 257.0551, 240.2677, 226.4221, 
      217.5795, 206.7036, 211.9852, 221.7744, 232.4703, 243.6246, 255.0728, 
      224.7775,
  227.4844, 205.5524, 223.0158, 244.1449, 241.3294, 230.7981, 224.0623, 
      220.5629, 218.7473, 218.6547, 221.0067, 227.8858, 239.3507, 252.4486, 
      186.8258 ;
  } // group GsiHofXBc

group: HofX {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  176.6368, 174.1857, 195.3052, 214.7622, 222.2356, 220.846, 216.4093, 
      213.2526, 209.9026, 207.9708, 208.2353, 212.4406, 220.8566, 233.73, 
      181.5446,
  166.8781, 159.7764, 224.5763, 255.6838, 252.8994, 238.6715, 227.2724, 
      218.4325, 212.0132, 215.4035, 221.0641, 228.2026, 237.0895, 246.2465, 
      223.784,
  292.9748, 293.4174, 286.41, 271.1309, 254.8238, 234.471, 220.8686, 
      210.5048, 204.9101, 213.452, 225.1687, 235.8813, 246.3493, 254.6549, 
      282.7286,
  153.0469, 155.6805, 220.744, 249.1663, 246.9592, 234.8852, 226.5111, 
      221.3778, 219.1345, 219.8379, 222.3798, 227.9497, 235.6271, 243.0406, 
      218.4219,
  275.6813, 274.0982, 277.9878, 272.5145, 261.0376, 242.5664, 228.1565, 
      215.6153, 203.5432, 209.8507, 221.3216, 233.3438, 243.8509, 253.2364, 
      283.7906,
  271.6429, 269.1485, 276.3429, 271.5592, 258.0934, 238.9886, 226.2866, 
      216.4929, 207.2805, 212.962, 223.3219, 233.0176, 240.6642, 247.7052, 
      284.5012,
  257.2548, 254.4906, 254.2988, 252.9041, 244.4244, 231.0509, 222.5009, 
      217.0181, 213.5159, 215.1574, 220.9328, 229.8975, 242.0261, 255.1175, 
      249.8248,
  185.7598, 171.108, 236.1643, 262.1205, 256.6778, 240.2876, 227.29, 
      216.6831, 207.5063, 212.584, 220.7504, 228.7155, 237.5468, 246.8313, 
      252.1144,
  267.3557, 268.3439, 268.8322, 261.2791, 249.7776, 233.4034, 222.6651, 
      215.5151, 212.2298, 215.4435, 222.5175, 231.7683, 241.7104, 251.5048, 
      267.7199,
  168.0432, 164.7606, 230.5948, 252.7646, 245.6549, 230.9738, 221.3597, 
      215.3269, 214.4045, 216.8591, 220.9403, 229.0795, 241.3861, 254.7864, 
      224.6138,
  158.0842, 164.4047, 224.3484, 246.5874, 244.68, 235.0927, 228.1079, 
      223.2104, 216.3487, 212.5453, 210.3054, 212.5406, 220.094, 232.3354, 
      228.6467,
  197.8513, 169.3049, 233.112, 264.0233, 259.5126, 242.1681, 227.9248, 
      215.7806, 204.4216, 210.5798, 221.9607, 234.3961, 246.1508, 256.0606, 
      250.1241,
  191.0477, 165.4345, 230.2722, 263.5005, 259.603, 242.2231, 227.8179, 
      215.5897, 203.9556, 209.6366, 221.415, 234.8128, 246.7379, 255.9029, 
      245.4932,
  182.6201, 165.8606, 230.6298, 258.8545, 253.7679, 237.7027, 225.6808, 
      216.6789, 210.7051, 215.2633, 224.1759, 234.5367, 245.0182, 255.5093, 
      238.6472,
  161.8278, 158.3778, 222.981, 251.5363, 249.4043, 236.8673, 227.0631, 
      219.7166, 213.1637, 213.8327, 217.3004, 223.9321, 233.2858, 243.4924, 
      226.0236,
  163.7971, 152.244, 219.926, 259.5825, 257.6855, 241.2264, 227.6269, 
      216.608, 207.0246, 212.0001, 221.7211, 232.1097, 242.7051, 253.7197, 
      220.5059,
  229.6282, 207.9446, 222.9126, 243.1598, 241.5118, 231.8967, 225.3438, 
      221.4922, 219.1168, 218.9814, 221.3634, 228.0966, 239.2607, 252.7536, 
      191.7876 ;
  } // group HofX

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -9223372036854775806LL ;
  		dateTime:units = "seconds since 2018-04-15T00:00:00Z" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  		string latitude:units = "degrees" ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  		string longitude:units = "degrees" ;
  	float sensorAzimuthAngle(Location) ;
  		sensorAzimuthAngle:_FillValue = 9.96921e+36f ;
  		string sensorAzimuthAngle:units = "degrees" ;
  	float sensorCentralFrequency(Channel) ;
  		sensorCentralFrequency:_FillValue = 9.96921e+36f ;
  		string sensorCentralFrequency:units = "Hz" ;
  	float sensorCentralWavenumber(Channel) ;
  		sensorCentralWavenumber:_FillValue = 9.96921e+36f ;
  		string sensorCentralWavenumber:units = "" ;
  	int sensorChannelNumber(Channel) ;
  		sensorChannelNumber:_FillValue = -2147483647 ;
  	int sensorPolarizationDirection(Channel) ;
  		sensorPolarizationDirection:_FillValue = -2147483647 ;
  	float sensorScanPosition(Location) ;
  		sensorScanPosition:_FillValue = 9.96921e+36f ;
  	float sensorViewAngle(Location) ;
  		sensorViewAngle:_FillValue = 9.96921e+36f ;
  		string sensorViewAngle:units = "degrees" ;
  	float sensorZenithAngle(Location) ;
  		sensorZenithAngle:_FillValue = 9.96921e+36f ;
  		string sensorZenithAngle:units = "degrees" ;
  	float solarAzimuthAngle(Location) ;
  		solarAzimuthAngle:_FillValue = 9.96921e+36f ;
  		string solarAzimuthAngle:units = "degrees" ;
  	float solarZenithAngle(Location) ;
  		solarZenithAngle:_FillValue = 9.96921e+36f ;
  		string solarZenithAngle:units = "degrees" ;
  data:

   dateTime = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16 ;

   latitude = -77.81, -42.5782, 12.6755, -47.5763, 4.7136, 26.5587, 60.6667, 
      -25.2042, 42.516, 50.4585, -63.0902, -9.7772, 0.5043, 26.6298, 
      -50.1559, -17.4598, 56.9285 ;

   longitude = 9.4296, 27.1671, 24.3545, 78.1395, 41.1401, 68.7682, 57.7598, 
      87.512, 82.3473, 200.5979, 227.6925, 208.5868, 234.0441, 202.8209, 
      247.2878, 261.8984, 266.1139 ;

   sensorAzimuthAngle = 296.67, 102.88, 281, 286.33, 96.05, 98.47, 105.47, 
      279.44, 286.06, 261.48, 72.55, 81.52, 260.26, 260.17, 78.92, 81.63, 
      250.46 ;

   sensorCentralFrequency = 23.79974, 31.4021, 50.30027, 52.80066, 53.59613, 
      54.40013, 54.93949, 55.49868, 57.29033, 57.29033, 57.29033, 57.29033, 
      57.29033, 57.29033, 89.01 ;

   sensorCentralWavenumber = 0.793874, 1.047461, 1.677836, 1.76124, 1.787774, 
      1.814593, 1.832584, 1.851237, 1.911, 1.911, 1.911, 1.911, 1.911, 1.911, 
      2.969054 ;

   sensorChannelNumber = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

   sensorPolarizationDirection = 9, 9, 9, 9, 10, 10, 9, 10, 10, 10, 10, 10, 
      10, 10, 9 ;

   sensorScanPosition = 8, 18, 4, 15, 16, 22, 19, 11, 8, 25, 13, 13, 18, 19, 
      15, 14, 16 ;

   sensorViewAngle = -25.002, 8.328, -38.334, -1.671, 1.662, 21.66, 11.661, 
      -15.003, -25.002, 31.659, -8.337, -8.337, 8.328, 11.661, -1.671, 
      -5.004, 1.662 ;

   sensorZenithAngle = -28.75, 9.48, -44.61, -1.89, 1.9, 24.72, 13.25, 
      -17.06, -28.6, 36.55, -9.5, -9.48, 9.46, 13.26, -1.9, -5.69, 1.89 ;

   solarAzimuthAngle = 144.79, 113.2, 74.73, 116.19, 76.12, 66.41, 69.46, 
      95.5, 70.71, 248.14, 288.32, 286.61, 280.89, 263.21, 292.12, 289.47, 
      234.58 ;

   solarZenithAngle = 109.79, 126.45, 109.58, 124.13, 119.33, 111.66, 90.24, 
      124.21, 96.32, 60.83, 91.69, 61.9, 60.08, 55.23, 84.6, 65.87, 58.54 ;
  } // group MetaData

group: ObsError {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5,
  2.5, 2.2, 2, 0.55, 0.3, 0.23, 0.23, 0.25, 0.25, 0.35, 0.4, 0.55, 0.8, 3, 
      3.5 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float brightnessTemperature(Location, Channel) ;
  		brightnessTemperature:_FillValue = 9.96921e+36f ;
  		string brightnessTemperature:units = "K" ;
  data:

   brightnessTemperature =
  172.21, 172.39, 193.94, 213.32, 219.62, 219.04, 215, 212.42, 208.86, 
      206.81, 207.34, 212.01, 221.1, 236.4, 181.98,
  175.54, 163.47, 227.25, 257.1, 253.83, 238, 225.91, 217.91, 210.3, 
      214.41, 220.74, 227.6, 236.86, 244.28, 229.08,
  276.32, 275.4, 274.81, 267.38, 252.57, 233.08, 218.67, 212.47, 203.51, 
      212.84, 224.06, 235.09, 245.57, 254.41, 271.36,
  147.09, 151.72, 217.65, 246.55, 245.6, 233.11, 224.51, 223.23, 218.97, 
      219.53, 222.41, 227.64, 235.62, 242.94, 210.6,
  278.3, 275.7, 278.7, 272.36, 260.37, 241.69, 226.91, 215.97, 202.77, 
      209.03, 220.71, 233.1, 244.68, 255.44, 283.76,
  284.81, 282.67, 282.51, 273.33, 258.1, 238.72, 225.44, 216.39, 205.62, 
      211.74, 222.81, 233.02, 240.48, 247.08, 286.51,
  256.61, 253.27, 253.59, 252.6, 243.78, 229.92, 221.87, 217.89, 212.94, 
      214.91, 221.05, 230.18, 243.1, 256.63, 247.65,
  169.99, 158.1, 225.58, 259.8, 256.13, 239.49, 226.63, 215.88, 207.21, 
      212.44, 220.95, 229.49, 238.2, 246.99, 227.76,
  243.62, 239.68, 243.81, 248.64, 244.18, 232.01, 221.67, 217.71, 211.48, 
      214.78, 222.61, 230.93, 242.97, 252.76, 235.42,
  165.92, 162.24, 228.42, 251.03, 244.53, 229.62, 219.98, 216.47, 213.33, 
      216.23, 219.8, 228.17, 241.47, 254.44, 221.38,
  152.71, 161.21, 219.46, 244.02, 243.31, 233.92, 227.1, 219.89, 216.86, 
      212.08, 209.54, 211.05, 218.78, 231.82, 213.86,
  203.27, 173.16, 235.41, 263.94, 258.87, 241.3, 227.53, 217.11, 203.65, 
      210.06, 221.3, 234.38, 246.22, 256.19, 253.71,
  193.64, 167.4, 231.78, 263.05, 258.77, 241.3, 226.13, 215.69, 202.54, 
      209.55, 221.41, 235.22, 247.29, 256.09, 247.56,
  186.81, 166.5, 230.39, 258.48, 253.71, 237.19, 224.99, 218.39, 210.04, 
      214.79, 223.99, 234.54, 244.34, 254.93, 237.76,
  173.44, 169.29, 231.43, 253.48, 249.6, 236.81, 225.83, 218.73, 211.66, 
      212.57, 216.62, 223.65, 232.4, 241.32, 244.47,
  161.29, 150.81, 218.88, 258.67, 256.95, 240.48, 226.22, 218.18, 206.96, 
      212.21, 222.19, 232.33, 243.77, 253.71, 216.83,
  235.57, 215.35, 230.25, 246.01, 241.71, 230.65, 225.22, 221.69, 218.46, 
      219.2, 221.24, 228.07, 239.01, 252.4, 198.56 ;
  } // group ObsValue
}
